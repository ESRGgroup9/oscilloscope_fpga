module Buffer2Pixel(
   input clk,
   input [7:0] R_i, G_i, B_i,

   output [23:0] pixel_o
);

endmodule

