// module top(

// );

// hdmiIP hdmiIP(
//    // clocks
//    .pixclk_i(pixclk_o),
//    .TMDS_clk_i(TMDS_clk_o),

//    .en_i(en_i),
//    .pixel_i(pixel_i),
//    // adc/filters output
//    .filteredSignal_i,

//    .TMDSp_o,
//    .TMDSn_o,
//    .TMDSp_clock_o,
//    .TMDSn_clock_o
// );